module main

import os

fn make_articles () []Article {
	mut articles := []Article{cap: 200}
	mut i := 1
	for fname in os.ls('data/') or { panic(err) }{
		articles << Article{
			id: i
			content: os.read_file('data/${fname}') or { panic(err) }
		}
		i += 1
	}
	return articles
}

fn make_articles2 () []Article{
	mut a := []Article{}
	a << Article{
		id: 1
		content: 'In an era where cyber attacks evolve faster than defenses, artificial intelligence is emerging as a game-changer in cybersecurity. Traditional antivirus software relies on signature-based detection, which struggles against zero-day exploits. AI, however, uses machine learning to analyze vast datasets in real-time, spotting anomalies like unusual network traffic or behavioral patterns indicative of malware.Consider a recent case where an AI system at a major bank flagged a sophisticated phishing attempt mid-transaction, preventing a multimillion-dollar loss. By training on historical breach data, AI predicts threats with up to 95% accuracy, far surpassing human analysts. Yet, challenges remain: AI models can be poisoned with adversarial inputs, leading to false positives or overlooked risks. As organizations integrate AI into security stacks, the key is hybrid approaches—combining human oversight with automated tools. The future? Proactive AI that not only detects but also autonomously neutralizes threats, reshaping digital fortresses worldwide.'
	}
	a << Article{
		id: 2
		content: "Quantum computers promise to revolutionize computation, but they pose a dire threat to current encryption standards. Algorithms like RSA and ECC, which secure online banking and communications, could be cracked in hours using Shor's algorithm on a sufficiently powerful quantum machine. Experts warn that harvest now, decrypt later attacks are already underway, with adversaries stockpiling encrypted data for future decryption. Governments are racing to develop post-quantum cryptography (PQC), with NIST standardizing algorithms like CRYSTALS-Kyber. Transitioning to PQC isn't simple—legacy systems must be audited, and key exchanges upgraded without disrupting services. While quantum tech is years away from breaking real-world encryption at scale, preparation is urgent. By 2030, experts predict widespread adoption of quantum-resistant protocols, ensuring data privacy endures the quantum leap."
	}
	a << Article{
		id: 3
		content: "The Internet of Things (IoT) connects billions of devices, from smart fridges to wearables, but convenience comes at a security cost. Many IoT gadgets ship with default passwords and unpatched firmware, turning them into easy entry points for hackers. A 2024 Mirai botnet variant hijacked over 500,000 unsecured cameras, launching DDoS attacks that crippled ISPs. Vulnerabilities often stem from rushed manufacturing—Chinese exports alone account for 70% of compromised devices due to lax standards. Mitigation starts with consumers: Change default credentials, enable two-factor authentication, and use network segmentation. On the industry side, regulations like the EU's Cyber Resilience Act mandate vulnerability disclosures. As IoT proliferates, robust security-by-design will be non-negotiable, preventing our connected homes from becoming hacker playgrounds."
	}
	a << Article{
		id: 4
		content: 'Ransomware has ballooned into a $20 billion industry, with groups like LockBit targeting hospitals and governments. Once crude encryptors, modern variants use double extortion—stealing data before locking it—forcing payouts via cryptocurrency. The 2025 Colonial Pipeline sequel hit a European energy firm, halting supplies for days. Attackers now employ living-off-the-land techniques, blending into legitimate tools to evade detection. Defenses are catching up: Endpoint detection platforms now incorporate behavioral analytics, while blockchain-based backups ensure immutable recovery. Governments are cracking down, with U.S. sanctions freezing ransomware wallets. The tide may turn as victim-sharing networks expose tactics, but until then, regular drills and zero-trust models remain essential shields against digital kidnappers.'
	}
	a << Article{
		id: 5
		content: 'Big data fuels innovation, from personalized ads to predictive healthcare, but it erodes privacy at an alarming rate. Companies like Meta harvest petabytes of user info, often without consent, enabling micro-targeted manipulation. The Cambridge Analytica scandal lingers as a cautionary tale, but 2025s breaches reveal deeper issues: AI-driven profiling infers sensitive details like political leanings from innocuous likes. GDPR fines have topped €2 billion, yet enforcement lags behind techs pace. Solutions include privacy-enhancing technologies (PETs) like homomorphic encryption, allowing data analysis without decryption. Users must demand transparency—opt for signal over noise in apps and support laws like Californias CCPA. In a world of constant data flows, reclaiming privacy means treating information as a fundamental right, not a commodity.'
	}
	a << Article{
		id: 6
		content: 'Blockchains immutable ledger, once synonymous with Bitcoin, is now fortifying global supply chains against fraud and tampering. By timestamping transactions across decentralized nodes, it ensures provenance—from farm to fork in food traceability. Walmarts IBM-partnered system reduced recall times from days to seconds during a 2024 E. coli outbreak, saving millions. In pharmaceuticals, blockchain verifies drug authenticity, combating counterfeit meds that kill 1 million annually. Challenges persist: Scalability limits throughput, and energy-intensive proof-of-work strains sustainability. Enterprise solutions like Hyperledger shift to permissioned networks for efficiency. As trade wars intensify, blockchains transparency could prevent disruptions, evolving from niche tech to a cornerstone of trustworthy commerce.'
	}
	a << Article{
		id: 7
		content: "5G's ultra-low latency promises transformative applications like autonomous vehicles, but its dense network architecture amplifies risks. With billions of new endpoints, the attack surface explodes—small cells become prime targets for signal jamming or man-in-the-middle intercepts. A simulated 2025 attack on a U.S. carrier demonstrated how rogue base stations could spoof towers, eavesdropping on calls. Spectrum sharing with military bands adds geopolitical tensions, as seen in Huawei bans. Security countermeasures include network slicing for isolated virtual networks and AI-monitored slicing for isolated virtual networks and AI-monitored traffic. Standards bodies like 3GPP are embedding zero-trust principles. As 5G blankets cities, balancing blistering speeds with ironclad defenses will define its legacy—innovation without isolation."
	}
	a << Article{
		id: 8
		content: 'Ethical hackers, or "white hats," are the unsung heroes probing systems for flaws before black hats exploit them. Bug bounty programs, like Google\'s, have paid out $50 million since 2010, uncovering vulnerabilities that could cost billions. In 2025, a teen hacker\'s report thwarted a nation-state cyber-espionage campaign targeting elections. Certifications like CEH train pros in penetration testing, simulating real attacks to harden defenses. Critics argue bounties incentivize chaos, but regulated platforms mitigate this. Governments now recruit ethical hackers for red-team exercises. As cyber threats democratize, empowering the good guys ensures a resilient digital ecosystem—turning potential breaches into fortified strengths.'
	}
	a << Article{
		id: 9
		content: 'Cloud adoption soars, with 94% of enterprises using multi-cloud setups, but misconfigurations cause 80% of breaches. Exposed S3 buckets in AWS have leaked sensitive data, from voter rolls to health records. Best practices emphasize shared responsibility: Providers secure infrastructure, but users must encrypt data at rest and enforce least-privilege access. Tools like AWS GuardDuty use ML to detect unauthorized API calls. The 2025 shift to confidential computing—processing encrypted data in trusted execution environments—promises ironclad privacy. For SMBs, managed services simplify compliance with standards like SOC 2. As clouds converge, proactive governance turns potential pitfalls into scalable sanctuaries.'
	}
	a << Article{
		id: 10
		content: 'Biometrics—fingerprints, face scans, iris patterns—are ditching passwords for seamless authentication, powering 70% of smartphones. Apple\'s Face ID uses 30,000+ infrared dots for spoof-proof recognition. Yet, deepfakes and 3D-printed masks challenge liveness detection, as a 2024 hack bypassed airport scanners. Privacy hawks decry centralized storage, vulnerable to breaches like the 2019 Suprema incident exposing 28 million fingerprints. Federated biometrics, storing templates on-device, mitigate risks, while multi-modal systems (face + voice) boost accuracy to 99.9%. Regulations like India\'s Aadhaar audits enforce ethical use. Biometrics herald a passwordless world, but only if we template trust with robust safeguards—securing identities without sacrificing souls.'
	}

	return a
}